/*****************************************************************************
 * ALU Flags
 * Copyright 2023 Anubhav Mattoo
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a
 * copy of this software and associated documentation files (the "Software"),
 * to deal in the Software without restriction, including without limitation
 * the rights to use, copy, modify, merge, publish, distribute, sublicense,
 * and/or sell copies of the Software, and to permit persons to whom the
 * Software is furnished to do so, subject to the following conditions:
 * 
 * The above copyright notice and this permission notice shall be included
 * in all copies or substantial portions of the Software.
 * 
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
 * FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
 * DEALINGS IN THE SOFTWARE.
 * 
 * Author : Anubhav Mattoo <anubhavmattoo@outlook.com>
 * Date : 2023 - 02 - 24
 ****************************************************************************/
 // `timescale 1ns/1ps


 module alu_flags (
	output [7:0] flags,
	 input [7:0] f,
	 input       a_b,
	 input       cn_n,
	 input       cn4_n,
	 input       cn8_n
);
	
	assign flags[0] = ~|f; // Zero
	assign flags[1] = ~cn8_n; // Carry
	assign flags[2] = a_b; // Equal
	assign flags[3] = ~cn_n & cn8_n; // Lesser Than
	assign flags[4] = cn_n & ~cn8_n; // Greater Than
	assign flags[5] = ~cn4_n; // Half Carry
	assign flags[6] = 0;
	assign flags[7] = 0;

endmodule